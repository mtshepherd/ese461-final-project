
module Top ( clk, reset, inputs, en, we, active_we, addr, wdata, output0, 
        output1, output2, output3, output4, output5, output6, output7, output8, 
        output9 );
  input [12543:0] inputs;
  input [1:0] en;
  input [793:0] we;
  input [17:0] addr;
  input [15:0] wdata;
  output [15:0] output0;
  output [15:0] output1;
  output [15:0] output2;
  output [15:0] output3;
  output [15:0] output4;
  output [15:0] output5;
  output [15:0] output6;
  output [15:0] output7;
  output [15:0] output8;
  output [15:0] output9;
  input clk, reset, active_we;
  wire   \l2[0].weights2[15] , \l2[0].weights2[14] , \l2[0].weights2[13] ,
         \l2[0].weights2[12] , \l2[0].weights2[11] , \l2[0].weights2[10] ,
         \l2[0].weights2[9] , \l2[0].weights2[8] , \l2[0].weights2[7] ,
         \l2[0].weights2[6] , \l2[0].weights2[5] , \l2[0].weights2[4] ,
         \l2[0].weights2[3] , \l2[0].weights2[2] , \l2[0].weights2[1] ,
         \l2[0].weights2[0] , \layer3pre[0][15] , \layer3pre[0][14] ,
         \layer3pre[0][13] , \layer3pre[0][12] , \layer3pre[0][11] ,
         \layer3pre[0][10] , \layer3pre[0][9] , \layer3pre[0][8] ,
         \layer3pre[0][7] , \layer3pre[0][6] , \layer3pre[0][5] ,
         \layer3pre[0][4] , \layer3pre[0][3] , \layer3pre[0][2] ,
         \layer3pre[0][1] , \layer3pre[0][0] , \layer3pre[1][15] ,
         \layer3pre[1][14] , \layer3pre[1][13] , \layer3pre[1][12] ,
         \layer3pre[1][11] , \layer3pre[1][10] , \layer3pre[1][9] ,
         \layer3pre[1][8] , \layer3pre[1][7] , \layer3pre[1][6] ,
         \layer3pre[1][5] , \layer3pre[1][4] , \layer3pre[1][3] ,
         \layer3pre[1][2] , \layer3pre[1][1] , \layer3pre[1][0] ,
         \layer3pre[2][15] , \layer3pre[2][14] , \layer3pre[2][13] ,
         \layer3pre[2][12] , \layer3pre[2][11] , \layer3pre[2][10] ,
         \layer3pre[2][9] , \layer3pre[2][8] , \layer3pre[2][7] ,
         \layer3pre[2][6] , \layer3pre[2][5] , \layer3pre[2][4] ,
         \layer3pre[2][3] , \layer3pre[2][2] , \layer3pre[2][1] ,
         \layer3pre[2][0] , \layer3pre[3][15] , \layer3pre[3][14] ,
         \layer3pre[3][13] , \layer3pre[3][12] , \layer3pre[3][11] ,
         \layer3pre[3][10] , \layer3pre[3][9] , \layer3pre[3][8] ,
         \layer3pre[3][7] , \layer3pre[3][6] , \layer3pre[3][5] ,
         \layer3pre[3][4] , \layer3pre[3][3] , \layer3pre[3][2] ,
         \layer3pre[3][1] , \layer3pre[3][0] , \layer3pre[4][15] ,
         \layer3pre[4][14] , \layer3pre[4][13] , \layer3pre[4][12] ,
         \layer3pre[4][11] , \layer3pre[4][10] , \layer3pre[4][9] ,
         \layer3pre[4][8] , \layer3pre[4][7] , \layer3pre[4][6] ,
         \layer3pre[4][5] , \layer3pre[4][4] , \layer3pre[4][3] ,
         \layer3pre[4][2] , \layer3pre[4][1] , \layer3pre[4][0] ,
         \layer3pre[5][15] , \layer3pre[5][14] , \layer3pre[5][13] ,
         \layer3pre[5][12] , \layer3pre[5][11] , \layer3pre[5][10] ,
         \layer3pre[5][9] , \layer3pre[5][8] , \layer3pre[5][7] ,
         \layer3pre[5][6] , \layer3pre[5][5] , \layer3pre[5][4] ,
         \layer3pre[5][3] , \layer3pre[5][2] , \layer3pre[5][1] ,
         \layer3pre[5][0] , \layer3pre[6][15] , \layer3pre[6][14] ,
         \layer3pre[6][13] , \layer3pre[6][12] , \layer3pre[6][11] ,
         \layer3pre[6][10] , \layer3pre[6][9] , \layer3pre[6][8] ,
         \layer3pre[6][7] , \layer3pre[6][6] , \layer3pre[6][5] ,
         \layer3pre[6][4] , \layer3pre[6][3] , \layer3pre[6][2] ,
         \layer3pre[6][1] , \layer3pre[6][0] , \layer3pre[7][15] ,
         \layer3pre[7][14] , \layer3pre[7][13] , \layer3pre[7][12] ,
         \layer3pre[7][11] , \layer3pre[7][10] , \layer3pre[7][9] ,
         \layer3pre[7][8] , \layer3pre[7][7] , \layer3pre[7][6] ,
         \layer3pre[7][5] , \layer3pre[7][4] , \layer3pre[7][3] ,
         \layer3pre[7][2] , \layer3pre[7][1] , \layer3pre[7][0] ,
         \layer3pre[8][15] , \layer3pre[8][14] , \layer3pre[8][13] ,
         \layer3pre[8][12] , \layer3pre[8][11] , \layer3pre[8][10] ,
         \layer3pre[8][9] , \layer3pre[8][8] , \layer3pre[8][7] ,
         \layer3pre[8][6] , \layer3pre[8][5] , \layer3pre[8][4] ,
         \layer3pre[8][3] , \layer3pre[8][2] , \layer3pre[8][1] ,
         \layer3pre[8][0] , \layer3pre[9][15] , \layer3pre[9][14] ,
         \layer3pre[9][13] , \layer3pre[9][12] , \layer3pre[9][11] ,
         \layer3pre[9][10] , \layer3pre[9][9] , \layer3pre[9][8] ,
         \layer3pre[9][7] , \layer3pre[9][6] , \layer3pre[9][5] ,
         \layer3pre[9][4] , \layer3pre[9][3] , \layer3pre[9][2] ,
         \layer3pre[9][1] , \layer3pre[9][0] , \l2[1].weights2[15] ,
         \l2[1].weights2[14] , \l2[1].weights2[13] , \l2[1].weights2[12] ,
         \l2[1].weights2[11] , \l2[1].weights2[10] , \l2[1].weights2[9] ,
         \l2[1].weights2[8] , \l2[1].weights2[7] , \l2[1].weights2[6] ,
         \l2[1].weights2[5] , \l2[1].weights2[4] , \l2[1].weights2[3] ,
         \l2[1].weights2[2] , \l2[1].weights2[1] , \l2[1].weights2[0] ,
         \l2[2].weights2[15] , \l2[2].weights2[14] , \l2[2].weights2[13] ,
         \l2[2].weights2[12] , \l2[2].weights2[11] , \l2[2].weights2[10] ,
         \l2[2].weights2[9] , \l2[2].weights2[8] , \l2[2].weights2[7] ,
         \l2[2].weights2[6] , \l2[2].weights2[5] , \l2[2].weights2[4] ,
         \l2[2].weights2[3] , \l2[2].weights2[2] , \l2[2].weights2[1] ,
         \l2[2].weights2[0] , \l2[3].weights2[15] , \l2[3].weights2[14] ,
         \l2[3].weights2[13] , \l2[3].weights2[12] , \l2[3].weights2[11] ,
         \l2[3].weights2[10] , \l2[3].weights2[9] , \l2[3].weights2[8] ,
         \l2[3].weights2[7] , \l2[3].weights2[6] , \l2[3].weights2[5] ,
         \l2[3].weights2[4] , \l2[3].weights2[3] , \l2[3].weights2[2] ,
         \l2[3].weights2[1] , \l2[3].weights2[0] , \l2[4].weights2[15] ,
         \l2[4].weights2[14] , \l2[4].weights2[13] , \l2[4].weights2[12] ,
         \l2[4].weights2[11] , \l2[4].weights2[10] , \l2[4].weights2[9] ,
         \l2[4].weights2[8] , \l2[4].weights2[7] , \l2[4].weights2[6] ,
         \l2[4].weights2[5] , \l2[4].weights2[4] , \l2[4].weights2[3] ,
         \l2[4].weights2[2] , \l2[4].weights2[1] , \l2[4].weights2[0] ,
         \l2[5].weights2[15] , \l2[5].weights2[14] , \l2[5].weights2[13] ,
         \l2[5].weights2[12] , \l2[5].weights2[11] , \l2[5].weights2[10] ,
         \l2[5].weights2[9] , \l2[5].weights2[8] , \l2[5].weights2[7] ,
         \l2[5].weights2[6] , \l2[5].weights2[5] , \l2[5].weights2[4] ,
         \l2[5].weights2[3] , \l2[5].weights2[2] , \l2[5].weights2[1] ,
         \l2[5].weights2[0] , \l2[6].weights2[15] , \l2[6].weights2[14] ,
         \l2[6].weights2[13] , \l2[6].weights2[12] , \l2[6].weights2[11] ,
         \l2[6].weights2[10] , \l2[6].weights2[9] , \l2[6].weights2[8] ,
         \l2[6].weights2[7] , \l2[6].weights2[6] , \l2[6].weights2[5] ,
         \l2[6].weights2[4] , \l2[6].weights2[3] , \l2[6].weights2[2] ,
         \l2[6].weights2[1] , \l2[6].weights2[0] , \l2[7].weights2[15] ,
         \l2[7].weights2[14] , \l2[7].weights2[13] , \l2[7].weights2[12] ,
         \l2[7].weights2[11] , \l2[7].weights2[10] , \l2[7].weights2[9] ,
         \l2[7].weights2[8] , \l2[7].weights2[7] , \l2[7].weights2[6] ,
         \l2[7].weights2[5] , \l2[7].weights2[4] , \l2[7].weights2[3] ,
         \l2[7].weights2[2] , \l2[7].weights2[1] , \l2[7].weights2[0] ,
         \l2[8].weights2[15] , \l2[8].weights2[14] , \l2[8].weights2[13] ,
         \l2[8].weights2[12] , \l2[8].weights2[11] , \l2[8].weights2[10] ,
         \l2[8].weights2[9] , \l2[8].weights2[8] , \l2[8].weights2[7] ,
         \l2[8].weights2[6] , \l2[8].weights2[5] , \l2[8].weights2[4] ,
         \l2[8].weights2[3] , \l2[8].weights2[2] , \l2[8].weights2[1] ,
         \l2[8].weights2[0] , \l2[9].weights2[15] , \l2[9].weights2[14] ,
         \l2[9].weights2[13] , \l2[9].weights2[12] , \l2[9].weights2[11] ,
         \l2[9].weights2[10] , \l2[9].weights2[9] , \l2[9].weights2[8] ,
         \l2[9].weights2[7] , \l2[9].weights2[6] , \l2[9].weights2[5] ,
         \l2[9].weights2[4] , \l2[9].weights2[3] , \l2[9].weights2[2] ,
         \l2[9].weights2[1] , \l2[9].weights2[0] ;
  wire   [15:0] layer1pre;
  wire   [15:0] layer1post;

  In_Calculator layer1 ( .p1(clk), .p2(reset), .p3(inputs), .p4(), .p5(
        layer1pre) );
  Activation active1 ( .p1(clk), .p2(active_we), .p3(layer1post), .p4(
        layer1pre), .p5(wdata) );
  ShiftRAM \l1[0].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[0]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[1].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[1]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[2].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[2]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[3].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[3]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[4].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[4]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[5].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[5]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[6].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[6]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[7].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[7]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[8].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[8]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[9].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[9]), 
        .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[10].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[10]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[11].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[11]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[12].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[12]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[13].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[13]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[14].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[14]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[15].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[15]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[16].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[16]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[17].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[17]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[18].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[18]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[19].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[19]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[20].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[20]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[21].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[21]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[22].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[22]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[23].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[23]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[24].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[24]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[25].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[25]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[26].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[26]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[27].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[27]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[28].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[28]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[29].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[29]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[30].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[30]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[31].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[31]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[32].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[32]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[33].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[33]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[34].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[34]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[35].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[35]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[36].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[36]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[37].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[37]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[38].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[38]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[39].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[39]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[40].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[40]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[41].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[41]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[42].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[42]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[43].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[43]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[44].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[44]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[45].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[45]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[46].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[46]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[47].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[47]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[48].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[48]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[49].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[49]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[50].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[50]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[51].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[51]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[52].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[52]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[53].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[53]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[54].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[54]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[55].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[55]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[56].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[56]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[57].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[57]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[58].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[58]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[59].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[59]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[60].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[60]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[61].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[61]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[62].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[62]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[63].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[63]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[64].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[64]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[65].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[65]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[66].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[66]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[67].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[67]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[68].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[68]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[69].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[69]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[70].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[70]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[71].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[71]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[72].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[72]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[73].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[73]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[74].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[74]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[75].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[75]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[76].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[76]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[77].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[77]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[78].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[78]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[79].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[79]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[80].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[80]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[81].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[81]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[82].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[82]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[83].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[83]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[84].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[84]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[85].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[85]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[86].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[86]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[87].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[87]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[88].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[88]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[89].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[89]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[90].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[90]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[91].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[91]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[92].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[92]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[93].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[93]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[94].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[94]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[95].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[95]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[96].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[96]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[97].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[97]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[98].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[98]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[99].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(we[99]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[100].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[100]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[101].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[101]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[102].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[102]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[103].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[103]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[104].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[104]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[105].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[105]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[106].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[106]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[107].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[107]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[108].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[108]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[109].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[109]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[110].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[110]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[111].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[111]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[112].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[112]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[113].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[113]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[114].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[114]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[115].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[115]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[116].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[116]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[117].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[117]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[118].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[118]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[119].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[119]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[120].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[120]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[121].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[121]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[122].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[122]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[123].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[123]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[124].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[124]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[125].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[125]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[126].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[126]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[127].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[127]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[128].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[128]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[129].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[129]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[130].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[130]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[131].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[131]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[132].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[132]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[133].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[133]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[134].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[134]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[135].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[135]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[136].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[136]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[137].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[137]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[138].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[138]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[139].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[139]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[140].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[140]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[141].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[141]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[142].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[142]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[143].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[143]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[144].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[144]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[145].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[145]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[146].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[146]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[147].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[147]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[148].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[148]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[149].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[149]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[150].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[150]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[151].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[151]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[152].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[152]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[153].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[153]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[154].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[154]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[155].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[155]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[156].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[156]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[157].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[157]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[158].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[158]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[159].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[159]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[160].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[160]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[161].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[161]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[162].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[162]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[163].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[163]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[164].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[164]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[165].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[165]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[166].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[166]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[167].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[167]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[168].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[168]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[169].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[169]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[170].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[170]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[171].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[171]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[172].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[172]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[173].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[173]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[174].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[174]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[175].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[175]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[176].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[176]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[177].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[177]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[178].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[178]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[179].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[179]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[180].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[180]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[181].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[181]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[182].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[182]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[183].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[183]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[184].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[184]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[185].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[185]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[186].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[186]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[187].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[187]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[188].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[188]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[189].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[189]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[190].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[190]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[191].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[191]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[192].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[192]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[193].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[193]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[194].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[194]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[195].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[195]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[196].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[196]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[197].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[197]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[198].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[198]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[199].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[199]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[200].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[200]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[201].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[201]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[202].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[202]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[203].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[203]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[204].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[204]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[205].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[205]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[206].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[206]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[207].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[207]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[208].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[208]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[209].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[209]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[210].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[210]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[211].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[211]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[212].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[212]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[213].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[213]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[214].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[214]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[215].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[215]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[216].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[216]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[217].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[217]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[218].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[218]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[219].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[219]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[220].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[220]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[221].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[221]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[222].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[222]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[223].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[223]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[224].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[224]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[225].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[225]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[226].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[226]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[227].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[227]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[228].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[228]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[229].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[229]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[230].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[230]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[231].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[231]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[232].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[232]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[233].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[233]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[234].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[234]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[235].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[235]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[236].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[236]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[237].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[237]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[238].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[238]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[239].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[239]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[240].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[240]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[241].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[241]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[242].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[242]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[243].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[243]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[244].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[244]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[245].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[245]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[246].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[246]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[247].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[247]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[248].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[248]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[249].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[249]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[250].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[250]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[251].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[251]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[252].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[252]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[253].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[253]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[254].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[254]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[255].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[255]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[256].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[256]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[257].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[257]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[258].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[258]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[259].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[259]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[260].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[260]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[261].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[261]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[262].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[262]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[263].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[263]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[264].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[264]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[265].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[265]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[266].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[266]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[267].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[267]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[268].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[268]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[269].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[269]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[270].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[270]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[271].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[271]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[272].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[272]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[273].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[273]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[274].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[274]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[275].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[275]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[276].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[276]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[277].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[277]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[278].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[278]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[279].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[279]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[280].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[280]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[281].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[281]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[282].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[282]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[283].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[283]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[284].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[284]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[285].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[285]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[286].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[286]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[287].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[287]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[288].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[288]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[289].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[289]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[290].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[290]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[291].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[291]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[292].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[292]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[293].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[293]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[294].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[294]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[295].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[295]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[296].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[296]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[297].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[297]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[298].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[298]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[299].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[299]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[300].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[300]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[301].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[301]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[302].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[302]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[303].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[303]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[304].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[304]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[305].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[305]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[306].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[306]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[307].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[307]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[308].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[308]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[309].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[309]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[310].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[310]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[311].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[311]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[312].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[312]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[313].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[313]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[314].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[314]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[315].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[315]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[316].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[316]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[317].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[317]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[318].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[318]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[319].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[319]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[320].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[320]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[321].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[321]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[322].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[322]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[323].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[323]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[324].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[324]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[325].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[325]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[326].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[326]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[327].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[327]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[328].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[328]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[329].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[329]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[330].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[330]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[331].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[331]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[332].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[332]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[333].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[333]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[334].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[334]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[335].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[335]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[336].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[336]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[337].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[337]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[338].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[338]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[339].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[339]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[340].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[340]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[341].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[341]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[342].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[342]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[343].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[343]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[344].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[344]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[345].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[345]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[346].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[346]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[347].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[347]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[348].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[348]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[349].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[349]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[350].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[350]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[351].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[351]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[352].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[352]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[353].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[353]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[354].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[354]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[355].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[355]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[356].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[356]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[357].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[357]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[358].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[358]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[359].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[359]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[360].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[360]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[361].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[361]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[362].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[362]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[363].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[363]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[364].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[364]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[365].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[365]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[366].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[366]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[367].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[367]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[368].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[368]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[369].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[369]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[370].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[370]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[371].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[371]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[372].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[372]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[373].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[373]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[374].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[374]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[375].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[375]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[376].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[376]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[377].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[377]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[378].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[378]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[379].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[379]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[380].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[380]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[381].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[381]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[382].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[382]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[383].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[383]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[384].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[384]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[385].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[385]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[386].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[386]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[387].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[387]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[388].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[388]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[389].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[389]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[390].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[390]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[391].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[391]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[392].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[392]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[393].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[393]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[394].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[394]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[395].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[395]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[396].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[396]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[397].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[397]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[398].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[398]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[399].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[399]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[400].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[400]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[401].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[401]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[402].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[402]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[403].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[403]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[404].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[404]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[405].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[405]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[406].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[406]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[407].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[407]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[408].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[408]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[409].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[409]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[410].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[410]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[411].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[411]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[412].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[412]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[413].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[413]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[414].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[414]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[415].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[415]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[416].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[416]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[417].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[417]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[418].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[418]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[419].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[419]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[420].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[420]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[421].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[421]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[422].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[422]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[423].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[423]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[424].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[424]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[425].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[425]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[426].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[426]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[427].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[427]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[428].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[428]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[429].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[429]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[430].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[430]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[431].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[431]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[432].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[432]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[433].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[433]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[434].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[434]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[435].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[435]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[436].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[436]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[437].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[437]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[438].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[438]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[439].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[439]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[440].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[440]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[441].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[441]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[442].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[442]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[443].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[443]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[444].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[444]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[445].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[445]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[446].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[446]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[447].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[447]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[448].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[448]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[449].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[449]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[450].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[450]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[451].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[451]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[452].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[452]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[453].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[453]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[454].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[454]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[455].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[455]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[456].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[456]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[457].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[457]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[458].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[458]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[459].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[459]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[460].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[460]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[461].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[461]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[462].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[462]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[463].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[463]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[464].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[464]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[465].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[465]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[466].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[466]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[467].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[467]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[468].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[468]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[469].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[469]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[470].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[470]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[471].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[471]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[472].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[472]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[473].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[473]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[474].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[474]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[475].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[475]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[476].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[476]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[477].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[477]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[478].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[478]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[479].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[479]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[480].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[480]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[481].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[481]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[482].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[482]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[483].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[483]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[484].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[484]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[485].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[485]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[486].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[486]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[487].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[487]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[488].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[488]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[489].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[489]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[490].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[490]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[491].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[491]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[492].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[492]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[493].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[493]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[494].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[494]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[495].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[495]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[496].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[496]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[497].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[497]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[498].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[498]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[499].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[499]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[500].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[500]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[501].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[501]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[502].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[502]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[503].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[503]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[504].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[504]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[505].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[505]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[506].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[506]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[507].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[507]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[508].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[508]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[509].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[509]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[510].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[510]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[511].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[511]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[512].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[512]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[513].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[513]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[514].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[514]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[515].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[515]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[516].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[516]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[517].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[517]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[518].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[518]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[519].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[519]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[520].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[520]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[521].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[521]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[522].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[522]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[523].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[523]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[524].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[524]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[525].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[525]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[526].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[526]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[527].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[527]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[528].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[528]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[529].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[529]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[530].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[530]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[531].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[531]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[532].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[532]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[533].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[533]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[534].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[534]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[535].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[535]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[536].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[536]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[537].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[537]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[538].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[538]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[539].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[539]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[540].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[540]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[541].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[541]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[542].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[542]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[543].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[543]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[544].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[544]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[545].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[545]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[546].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[546]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[547].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[547]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[548].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[548]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[549].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[549]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[550].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[550]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[551].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[551]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[552].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[552]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[553].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[553]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[554].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[554]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[555].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[555]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[556].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[556]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[557].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[557]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[558].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[558]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[559].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[559]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[560].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[560]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[561].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[561]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[562].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[562]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[563].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[563]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[564].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[564]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[565].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[565]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[566].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[566]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[567].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[567]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[568].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[568]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[569].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[569]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[570].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[570]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[571].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[571]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[572].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[572]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[573].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[573]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[574].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[574]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[575].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[575]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[576].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[576]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[577].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[577]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[578].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[578]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[579].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[579]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[580].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[580]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[581].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[581]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[582].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[582]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[583].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[583]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[584].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[584]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[585].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[585]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[586].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[586]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[587].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[587]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[588].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[588]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[589].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[589]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[590].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[590]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[591].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[591]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[592].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[592]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[593].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[593]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[594].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[594]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[595].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[595]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[596].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[596]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[597].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[597]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[598].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[598]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[599].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[599]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[600].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[600]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[601].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[601]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[602].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[602]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[603].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[603]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[604].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[604]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[605].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[605]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[606].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[606]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[607].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[607]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[608].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[608]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[609].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[609]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[610].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[610]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[611].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[611]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[612].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[612]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[613].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[613]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[614].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[614]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[615].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[615]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[616].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[616]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[617].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[617]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[618].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[618]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[619].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[619]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[620].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[620]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[621].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[621]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[622].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[622]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[623].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[623]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[624].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[624]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[625].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[625]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[626].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[626]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[627].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[627]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[628].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[628]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[629].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[629]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[630].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[630]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[631].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[631]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[632].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[632]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[633].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[633]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[634].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[634]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[635].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[635]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[636].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[636]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[637].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[637]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[638].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[638]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[639].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[639]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[640].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[640]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[641].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[641]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[642].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[642]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[643].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[643]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[644].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[644]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[645].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[645]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[646].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[646]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[647].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[647]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[648].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[648]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[649].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[649]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[650].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[650]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[651].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[651]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[652].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[652]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[653].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[653]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[654].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[654]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[655].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[655]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[656].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[656]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[657].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[657]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[658].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[658]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[659].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[659]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[660].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[660]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[661].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[661]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[662].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[662]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[663].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[663]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[664].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[664]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[665].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[665]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[666].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[666]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[667].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[667]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[668].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[668]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[669].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[669]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[670].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[670]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[671].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[671]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[672].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[672]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[673].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[673]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[674].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[674]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[675].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[675]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[676].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[676]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[677].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[677]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[678].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[678]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[679].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[679]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[680].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[680]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[681].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[681]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[682].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[682]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[683].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[683]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[684].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[684]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[685].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[685]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[686].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[686]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[687].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[687]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[688].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[688]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[689].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[689]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[690].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[690]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[691].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[691]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[692].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[692]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[693].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[693]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[694].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[694]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[695].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[695]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[696].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[696]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[697].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[697]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[698].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[698]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[699].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[699]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[700].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[700]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[701].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[701]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[702].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[702]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[703].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[703]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[704].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[704]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[705].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[705]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[706].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[706]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[707].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[707]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[708].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[708]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[709].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[709]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[710].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[710]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[711].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[711]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[712].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[712]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[713].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[713]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[714].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[714]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[715].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[715]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[716].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[716]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[717].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[717]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[718].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[718]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[719].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[719]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[720].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[720]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[721].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[721]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[722].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[722]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[723].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[723]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[724].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[724]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[725].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[725]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[726].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[726]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[727].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[727]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[728].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[728]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[729].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[729]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[730].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[730]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[731].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[731]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[732].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[732]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[733].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[733]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[734].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[734]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[735].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[735]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[736].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[736]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[737].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[737]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[738].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[738]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[739].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[739]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[740].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[740]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[741].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[741]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[742].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[742]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[743].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[743]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[744].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[744]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[745].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[745]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[746].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[746]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[747].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[747]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[748].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[748]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[749].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[749]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[750].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[750]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[751].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[751]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[752].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[752]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[753].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[753]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[754].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[754]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[755].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[755]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[756].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[756]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[757].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[757]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[758].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[758]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[759].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[759]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[760].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[760]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[761].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[761]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[762].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[762]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[763].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[763]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[764].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[764]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[765].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[765]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[766].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[766]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[767].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[767]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[768].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[768]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[769].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[769]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[770].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[770]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[771].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[771]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[772].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[772]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[773].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[773]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[774].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[774]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[775].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[775]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[776].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[776]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[777].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[777]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[778].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[778]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[779].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[779]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[780].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[780]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[781].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[781]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[782].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[782]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l1[783].weightsRAM1  ( .p1(clk), .p2(reset), .p3(en[0]), .p4(
        we[783]), .p5(), .p6(addr), .p7(wdata) );
  ShiftRAM \l2[0].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[784]), .p5({\l2[0].weights2[15] , \l2[0].weights2[14] , \l2[0].weights2[13] , 
        \l2[0].weights2[12] , \l2[0].weights2[11] , \l2[0].weights2[10] , 
        \l2[0].weights2[9] , \l2[0].weights2[8] , \l2[0].weights2[7] , 
        \l2[0].weights2[6] , \l2[0].weights2[5] , \l2[0].weights2[4] , 
        \l2[0].weights2[3] , \l2[0].weights2[2] , \l2[0].weights2[1] , 
        \l2[0].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[0].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[0].weights2[15] , \l2[0].weights2[14] , \l2[0].weights2[13] , 
        \l2[0].weights2[12] , \l2[0].weights2[11] , \l2[0].weights2[10] , 
        \l2[0].weights2[9] , \l2[0].weights2[8] , \l2[0].weights2[7] , 
        \l2[0].weights2[6] , \l2[0].weights2[5] , \l2[0].weights2[4] , 
        \l2[0].weights2[3] , \l2[0].weights2[2] , \l2[0].weights2[1] , 
        \l2[0].weights2[0] }), .p5({\layer3pre[0][15] , \layer3pre[0][14] , 
        \layer3pre[0][13] , \layer3pre[0][12] , \layer3pre[0][11] , 
        \layer3pre[0][10] , \layer3pre[0][9] , \layer3pre[0][8] , 
        \layer3pre[0][7] , \layer3pre[0][6] , \layer3pre[0][5] , 
        \layer3pre[0][4] , \layer3pre[0][3] , \layer3pre[0][2] , 
        \layer3pre[0][1] , \layer3pre[0][0] }) );
  Activation \l2[0].active2  ( .p1(clk), .p2(active_we), .p3(output0), .p4({
        \layer3pre[0][15] , \layer3pre[0][14] , \layer3pre[0][13] , 
        \layer3pre[0][12] , \layer3pre[0][11] , \layer3pre[0][10] , 
        \layer3pre[0][9] , \layer3pre[0][8] , \layer3pre[0][7] , 
        \layer3pre[0][6] , \layer3pre[0][5] , \layer3pre[0][4] , 
        \layer3pre[0][3] , \layer3pre[0][2] , \layer3pre[0][1] , 
        \layer3pre[0][0] }), .p5(wdata) );
  ShiftRAM \l2[1].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[785]), .p5({\l2[1].weights2[15] , \l2[1].weights2[14] , \l2[1].weights2[13] , 
        \l2[1].weights2[12] , \l2[1].weights2[11] , \l2[1].weights2[10] , 
        \l2[1].weights2[9] , \l2[1].weights2[8] , \l2[1].weights2[7] , 
        \l2[1].weights2[6] , \l2[1].weights2[5] , \l2[1].weights2[4] , 
        \l2[1].weights2[3] , \l2[1].weights2[2] , \l2[1].weights2[1] , 
        \l2[1].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[1].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[1].weights2[15] , \l2[1].weights2[14] , \l2[1].weights2[13] , 
        \l2[1].weights2[12] , \l2[1].weights2[11] , \l2[1].weights2[10] , 
        \l2[1].weights2[9] , \l2[1].weights2[8] , \l2[1].weights2[7] , 
        \l2[1].weights2[6] , \l2[1].weights2[5] , \l2[1].weights2[4] , 
        \l2[1].weights2[3] , \l2[1].weights2[2] , \l2[1].weights2[1] , 
        \l2[1].weights2[0] }), .p5({\layer3pre[1][15] , \layer3pre[1][14] , 
        \layer3pre[1][13] , \layer3pre[1][12] , \layer3pre[1][11] , 
        \layer3pre[1][10] , \layer3pre[1][9] , \layer3pre[1][8] , 
        \layer3pre[1][7] , \layer3pre[1][6] , \layer3pre[1][5] , 
        \layer3pre[1][4] , \layer3pre[1][3] , \layer3pre[1][2] , 
        \layer3pre[1][1] , \layer3pre[1][0] }) );
  Activation \l2[1].active2  ( .p1(clk), .p2(active_we), .p3(output1), .p4({
        \layer3pre[1][15] , \layer3pre[1][14] , \layer3pre[1][13] , 
        \layer3pre[1][12] , \layer3pre[1][11] , \layer3pre[1][10] , 
        \layer3pre[1][9] , \layer3pre[1][8] , \layer3pre[1][7] , 
        \layer3pre[1][6] , \layer3pre[1][5] , \layer3pre[1][4] , 
        \layer3pre[1][3] , \layer3pre[1][2] , \layer3pre[1][1] , 
        \layer3pre[1][0] }), .p5(wdata) );
  ShiftRAM \l2[2].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[786]), .p5({\l2[2].weights2[15] , \l2[2].weights2[14] , \l2[2].weights2[13] , 
        \l2[2].weights2[12] , \l2[2].weights2[11] , \l2[2].weights2[10] , 
        \l2[2].weights2[9] , \l2[2].weights2[8] , \l2[2].weights2[7] , 
        \l2[2].weights2[6] , \l2[2].weights2[5] , \l2[2].weights2[4] , 
        \l2[2].weights2[3] , \l2[2].weights2[2] , \l2[2].weights2[1] , 
        \l2[2].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[2].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[2].weights2[15] , \l2[2].weights2[14] , \l2[2].weights2[13] , 
        \l2[2].weights2[12] , \l2[2].weights2[11] , \l2[2].weights2[10] , 
        \l2[2].weights2[9] , \l2[2].weights2[8] , \l2[2].weights2[7] , 
        \l2[2].weights2[6] , \l2[2].weights2[5] , \l2[2].weights2[4] , 
        \l2[2].weights2[3] , \l2[2].weights2[2] , \l2[2].weights2[1] , 
        \l2[2].weights2[0] }), .p5({\layer3pre[2][15] , \layer3pre[2][14] , 
        \layer3pre[2][13] , \layer3pre[2][12] , \layer3pre[2][11] , 
        \layer3pre[2][10] , \layer3pre[2][9] , \layer3pre[2][8] , 
        \layer3pre[2][7] , \layer3pre[2][6] , \layer3pre[2][5] , 
        \layer3pre[2][4] , \layer3pre[2][3] , \layer3pre[2][2] , 
        \layer3pre[2][1] , \layer3pre[2][0] }) );
  Activation \l2[2].active2  ( .p1(clk), .p2(active_we), .p3(output2), .p4({
        \layer3pre[2][15] , \layer3pre[2][14] , \layer3pre[2][13] , 
        \layer3pre[2][12] , \layer3pre[2][11] , \layer3pre[2][10] , 
        \layer3pre[2][9] , \layer3pre[2][8] , \layer3pre[2][7] , 
        \layer3pre[2][6] , \layer3pre[2][5] , \layer3pre[2][4] , 
        \layer3pre[2][3] , \layer3pre[2][2] , \layer3pre[2][1] , 
        \layer3pre[2][0] }), .p5(wdata) );
  ShiftRAM \l2[3].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[787]), .p5({\l2[3].weights2[15] , \l2[3].weights2[14] , \l2[3].weights2[13] , 
        \l2[3].weights2[12] , \l2[3].weights2[11] , \l2[3].weights2[10] , 
        \l2[3].weights2[9] , \l2[3].weights2[8] , \l2[3].weights2[7] , 
        \l2[3].weights2[6] , \l2[3].weights2[5] , \l2[3].weights2[4] , 
        \l2[3].weights2[3] , \l2[3].weights2[2] , \l2[3].weights2[1] , 
        \l2[3].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[3].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[3].weights2[15] , \l2[3].weights2[14] , \l2[3].weights2[13] , 
        \l2[3].weights2[12] , \l2[3].weights2[11] , \l2[3].weights2[10] , 
        \l2[3].weights2[9] , \l2[3].weights2[8] , \l2[3].weights2[7] , 
        \l2[3].weights2[6] , \l2[3].weights2[5] , \l2[3].weights2[4] , 
        \l2[3].weights2[3] , \l2[3].weights2[2] , \l2[3].weights2[1] , 
        \l2[3].weights2[0] }), .p5({\layer3pre[3][15] , \layer3pre[3][14] , 
        \layer3pre[3][13] , \layer3pre[3][12] , \layer3pre[3][11] , 
        \layer3pre[3][10] , \layer3pre[3][9] , \layer3pre[3][8] , 
        \layer3pre[3][7] , \layer3pre[3][6] , \layer3pre[3][5] , 
        \layer3pre[3][4] , \layer3pre[3][3] , \layer3pre[3][2] , 
        \layer3pre[3][1] , \layer3pre[3][0] }) );
  Activation \l2[3].active2  ( .p1(clk), .p2(active_we), .p3(output3), .p4({
        \layer3pre[3][15] , \layer3pre[3][14] , \layer3pre[3][13] , 
        \layer3pre[3][12] , \layer3pre[3][11] , \layer3pre[3][10] , 
        \layer3pre[3][9] , \layer3pre[3][8] , \layer3pre[3][7] , 
        \layer3pre[3][6] , \layer3pre[3][5] , \layer3pre[3][4] , 
        \layer3pre[3][3] , \layer3pre[3][2] , \layer3pre[3][1] , 
        \layer3pre[3][0] }), .p5(wdata) );
  ShiftRAM \l2[4].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[788]), .p5({\l2[4].weights2[15] , \l2[4].weights2[14] , \l2[4].weights2[13] , 
        \l2[4].weights2[12] , \l2[4].weights2[11] , \l2[4].weights2[10] , 
        \l2[4].weights2[9] , \l2[4].weights2[8] , \l2[4].weights2[7] , 
        \l2[4].weights2[6] , \l2[4].weights2[5] , \l2[4].weights2[4] , 
        \l2[4].weights2[3] , \l2[4].weights2[2] , \l2[4].weights2[1] , 
        \l2[4].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[4].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[4].weights2[15] , \l2[4].weights2[14] , \l2[4].weights2[13] , 
        \l2[4].weights2[12] , \l2[4].weights2[11] , \l2[4].weights2[10] , 
        \l2[4].weights2[9] , \l2[4].weights2[8] , \l2[4].weights2[7] , 
        \l2[4].weights2[6] , \l2[4].weights2[5] , \l2[4].weights2[4] , 
        \l2[4].weights2[3] , \l2[4].weights2[2] , \l2[4].weights2[1] , 
        \l2[4].weights2[0] }), .p5({\layer3pre[4][15] , \layer3pre[4][14] , 
        \layer3pre[4][13] , \layer3pre[4][12] , \layer3pre[4][11] , 
        \layer3pre[4][10] , \layer3pre[4][9] , \layer3pre[4][8] , 
        \layer3pre[4][7] , \layer3pre[4][6] , \layer3pre[4][5] , 
        \layer3pre[4][4] , \layer3pre[4][3] , \layer3pre[4][2] , 
        \layer3pre[4][1] , \layer3pre[4][0] }) );
  Activation \l2[4].active2  ( .p1(clk), .p2(active_we), .p3(output4), .p4({
        \layer3pre[4][15] , \layer3pre[4][14] , \layer3pre[4][13] , 
        \layer3pre[4][12] , \layer3pre[4][11] , \layer3pre[4][10] , 
        \layer3pre[4][9] , \layer3pre[4][8] , \layer3pre[4][7] , 
        \layer3pre[4][6] , \layer3pre[4][5] , \layer3pre[4][4] , 
        \layer3pre[4][3] , \layer3pre[4][2] , \layer3pre[4][1] , 
        \layer3pre[4][0] }), .p5(wdata) );
  ShiftRAM \l2[5].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[789]), .p5({\l2[5].weights2[15] , \l2[5].weights2[14] , \l2[5].weights2[13] , 
        \l2[5].weights2[12] , \l2[5].weights2[11] , \l2[5].weights2[10] , 
        \l2[5].weights2[9] , \l2[5].weights2[8] , \l2[5].weights2[7] , 
        \l2[5].weights2[6] , \l2[5].weights2[5] , \l2[5].weights2[4] , 
        \l2[5].weights2[3] , \l2[5].weights2[2] , \l2[5].weights2[1] , 
        \l2[5].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[5].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[5].weights2[15] , \l2[5].weights2[14] , \l2[5].weights2[13] , 
        \l2[5].weights2[12] , \l2[5].weights2[11] , \l2[5].weights2[10] , 
        \l2[5].weights2[9] , \l2[5].weights2[8] , \l2[5].weights2[7] , 
        \l2[5].weights2[6] , \l2[5].weights2[5] , \l2[5].weights2[4] , 
        \l2[5].weights2[3] , \l2[5].weights2[2] , \l2[5].weights2[1] , 
        \l2[5].weights2[0] }), .p5({\layer3pre[5][15] , \layer3pre[5][14] , 
        \layer3pre[5][13] , \layer3pre[5][12] , \layer3pre[5][11] , 
        \layer3pre[5][10] , \layer3pre[5][9] , \layer3pre[5][8] , 
        \layer3pre[5][7] , \layer3pre[5][6] , \layer3pre[5][5] , 
        \layer3pre[5][4] , \layer3pre[5][3] , \layer3pre[5][2] , 
        \layer3pre[5][1] , \layer3pre[5][0] }) );
  Activation \l2[5].active2  ( .p1(clk), .p2(active_we), .p3(output5), .p4({
        \layer3pre[5][15] , \layer3pre[5][14] , \layer3pre[5][13] , 
        \layer3pre[5][12] , \layer3pre[5][11] , \layer3pre[5][10] , 
        \layer3pre[5][9] , \layer3pre[5][8] , \layer3pre[5][7] , 
        \layer3pre[5][6] , \layer3pre[5][5] , \layer3pre[5][4] , 
        \layer3pre[5][3] , \layer3pre[5][2] , \layer3pre[5][1] , 
        \layer3pre[5][0] }), .p5(wdata) );
  ShiftRAM \l2[6].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[790]), .p5({\l2[6].weights2[15] , \l2[6].weights2[14] , \l2[6].weights2[13] , 
        \l2[6].weights2[12] , \l2[6].weights2[11] , \l2[6].weights2[10] , 
        \l2[6].weights2[9] , \l2[6].weights2[8] , \l2[6].weights2[7] , 
        \l2[6].weights2[6] , \l2[6].weights2[5] , \l2[6].weights2[4] , 
        \l2[6].weights2[3] , \l2[6].weights2[2] , \l2[6].weights2[1] , 
        \l2[6].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[6].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[6].weights2[15] , \l2[6].weights2[14] , \l2[6].weights2[13] , 
        \l2[6].weights2[12] , \l2[6].weights2[11] , \l2[6].weights2[10] , 
        \l2[6].weights2[9] , \l2[6].weights2[8] , \l2[6].weights2[7] , 
        \l2[6].weights2[6] , \l2[6].weights2[5] , \l2[6].weights2[4] , 
        \l2[6].weights2[3] , \l2[6].weights2[2] , \l2[6].weights2[1] , 
        \l2[6].weights2[0] }), .p5({\layer3pre[6][15] , \layer3pre[6][14] , 
        \layer3pre[6][13] , \layer3pre[6][12] , \layer3pre[6][11] , 
        \layer3pre[6][10] , \layer3pre[6][9] , \layer3pre[6][8] , 
        \layer3pre[6][7] , \layer3pre[6][6] , \layer3pre[6][5] , 
        \layer3pre[6][4] , \layer3pre[6][3] , \layer3pre[6][2] , 
        \layer3pre[6][1] , \layer3pre[6][0] }) );
  Activation \l2[6].active2  ( .p1(clk), .p2(active_we), .p3(output6), .p4({
        \layer3pre[6][15] , \layer3pre[6][14] , \layer3pre[6][13] , 
        \layer3pre[6][12] , \layer3pre[6][11] , \layer3pre[6][10] , 
        \layer3pre[6][9] , \layer3pre[6][8] , \layer3pre[6][7] , 
        \layer3pre[6][6] , \layer3pre[6][5] , \layer3pre[6][4] , 
        \layer3pre[6][3] , \layer3pre[6][2] , \layer3pre[6][1] , 
        \layer3pre[6][0] }), .p5(wdata) );
  ShiftRAM \l2[7].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[791]), .p5({\l2[7].weights2[15] , \l2[7].weights2[14] , \l2[7].weights2[13] , 
        \l2[7].weights2[12] , \l2[7].weights2[11] , \l2[7].weights2[10] , 
        \l2[7].weights2[9] , \l2[7].weights2[8] , \l2[7].weights2[7] , 
        \l2[7].weights2[6] , \l2[7].weights2[5] , \l2[7].weights2[4] , 
        \l2[7].weights2[3] , \l2[7].weights2[2] , \l2[7].weights2[1] , 
        \l2[7].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[7].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[7].weights2[15] , \l2[7].weights2[14] , \l2[7].weights2[13] , 
        \l2[7].weights2[12] , \l2[7].weights2[11] , \l2[7].weights2[10] , 
        \l2[7].weights2[9] , \l2[7].weights2[8] , \l2[7].weights2[7] , 
        \l2[7].weights2[6] , \l2[7].weights2[5] , \l2[7].weights2[4] , 
        \l2[7].weights2[3] , \l2[7].weights2[2] , \l2[7].weights2[1] , 
        \l2[7].weights2[0] }), .p5({\layer3pre[7][15] , \layer3pre[7][14] , 
        \layer3pre[7][13] , \layer3pre[7][12] , \layer3pre[7][11] , 
        \layer3pre[7][10] , \layer3pre[7][9] , \layer3pre[7][8] , 
        \layer3pre[7][7] , \layer3pre[7][6] , \layer3pre[7][5] , 
        \layer3pre[7][4] , \layer3pre[7][3] , \layer3pre[7][2] , 
        \layer3pre[7][1] , \layer3pre[7][0] }) );
  Activation \l2[7].active2  ( .p1(clk), .p2(active_we), .p3(output7), .p4({
        \layer3pre[7][15] , \layer3pre[7][14] , \layer3pre[7][13] , 
        \layer3pre[7][12] , \layer3pre[7][11] , \layer3pre[7][10] , 
        \layer3pre[7][9] , \layer3pre[7][8] , \layer3pre[7][7] , 
        \layer3pre[7][6] , \layer3pre[7][5] , \layer3pre[7][4] , 
        \layer3pre[7][3] , \layer3pre[7][2] , \layer3pre[7][1] , 
        \layer3pre[7][0] }), .p5(wdata) );
  ShiftRAM \l2[8].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[792]), .p5({\l2[8].weights2[15] , \l2[8].weights2[14] , \l2[8].weights2[13] , 
        \l2[8].weights2[12] , \l2[8].weights2[11] , \l2[8].weights2[10] , 
        \l2[8].weights2[9] , \l2[8].weights2[8] , \l2[8].weights2[7] , 
        \l2[8].weights2[6] , \l2[8].weights2[5] , \l2[8].weights2[4] , 
        \l2[8].weights2[3] , \l2[8].weights2[2] , \l2[8].weights2[1] , 
        \l2[8].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[8].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[8].weights2[15] , \l2[8].weights2[14] , \l2[8].weights2[13] , 
        \l2[8].weights2[12] , \l2[8].weights2[11] , \l2[8].weights2[10] , 
        \l2[8].weights2[9] , \l2[8].weights2[8] , \l2[8].weights2[7] , 
        \l2[8].weights2[6] , \l2[8].weights2[5] , \l2[8].weights2[4] , 
        \l2[8].weights2[3] , \l2[8].weights2[2] , \l2[8].weights2[1] , 
        \l2[8].weights2[0] }), .p5({\layer3pre[8][15] , \layer3pre[8][14] , 
        \layer3pre[8][13] , \layer3pre[8][12] , \layer3pre[8][11] , 
        \layer3pre[8][10] , \layer3pre[8][9] , \layer3pre[8][8] , 
        \layer3pre[8][7] , \layer3pre[8][6] , \layer3pre[8][5] , 
        \layer3pre[8][4] , \layer3pre[8][3] , \layer3pre[8][2] , 
        \layer3pre[8][1] , \layer3pre[8][0] }) );
  Activation \l2[8].active2  ( .p1(clk), .p2(active_we), .p3(output8), .p4({
        \layer3pre[8][15] , \layer3pre[8][14] , \layer3pre[8][13] , 
        \layer3pre[8][12] , \layer3pre[8][11] , \layer3pre[8][10] , 
        \layer3pre[8][9] , \layer3pre[8][8] , \layer3pre[8][7] , 
        \layer3pre[8][6] , \layer3pre[8][5] , \layer3pre[8][4] , 
        \layer3pre[8][3] , \layer3pre[8][2] , \layer3pre[8][1] , 
        \layer3pre[8][0] }), .p5(wdata) );
  ShiftRAM \l2[9].weightsRAM2  ( .p1(clk), .p2(reset), .p3(en[1]), .p4(we[793]), .p5({\l2[9].weights2[15] , \l2[9].weights2[14] , \l2[9].weights2[13] , 
        \l2[9].weights2[12] , \l2[9].weights2[11] , \l2[9].weights2[10] , 
        \l2[9].weights2[9] , \l2[9].weights2[8] , \l2[9].weights2[7] , 
        \l2[9].weights2[6] , \l2[9].weights2[5] , \l2[9].weights2[4] , 
        \l2[9].weights2[3] , \l2[9].weights2[2] , \l2[9].weights2[1] , 
        \l2[9].weights2[0] }), .p6(addr), .p7(wdata) );
  Out_Calculator \l2[9].layer2  ( .p1(clk), .p2(reset), .p3(layer1post), .p4({
        \l2[9].weights2[15] , \l2[9].weights2[14] , \l2[9].weights2[13] , 
        \l2[9].weights2[12] , \l2[9].weights2[11] , \l2[9].weights2[10] , 
        \l2[9].weights2[9] , \l2[9].weights2[8] , \l2[9].weights2[7] , 
        \l2[9].weights2[6] , \l2[9].weights2[5] , \l2[9].weights2[4] , 
        \l2[9].weights2[3] , \l2[9].weights2[2] , \l2[9].weights2[1] , 
        \l2[9].weights2[0] }), .p5({\layer3pre[9][15] , \layer3pre[9][14] , 
        \layer3pre[9][13] , \layer3pre[9][12] , \layer3pre[9][11] , 
        \layer3pre[9][10] , \layer3pre[9][9] , \layer3pre[9][8] , 
        \layer3pre[9][7] , \layer3pre[9][6] , \layer3pre[9][5] , 
        \layer3pre[9][4] , \layer3pre[9][3] , \layer3pre[9][2] , 
        \layer3pre[9][1] , \layer3pre[9][0] }) );
  Activation \l2[9].active2  ( .p1(clk), .p2(active_we), .p3(output9), .p4({
        \layer3pre[9][15] , \layer3pre[9][14] , \layer3pre[9][13] , 
        \layer3pre[9][12] , \layer3pre[9][11] , \layer3pre[9][10] , 
        \layer3pre[9][9] , \layer3pre[9][8] , \layer3pre[9][7] , 
        \layer3pre[9][6] , \layer3pre[9][5] , \layer3pre[9][4] , 
        \layer3pre[9][3] , \layer3pre[9][2] , \layer3pre[9][1] , 
        \layer3pre[9][0] }), .p5(wdata) );
endmodule

